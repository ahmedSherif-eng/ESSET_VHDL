library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity ConditionalByPass is
    generic (
        OUTPUT_SIZE : integer := 8  -- Default output size is 32 bits
    );
    port (
        clk       : in  std_logic;
        i_DV      : in  std_logic;
        o_status  : out std_logic; -- condition found or not
        i_input   : in  std_logic_vector(OUTPUT_SIZE - 1 downto 0)
    );
end ConditionalByPass;

architecture behav of ConditionalByPass is
    signal r_input     : std_logic_vector(OUTPUT_SIZE - 1 downto 0) := (others => '0');
    signal r_condition : std_logic_vector(OUTPUT_SIZE - 1 downto 0) := X"33";
    signal r_status    : std_logic := '0';
    --signal r_first     : std_logic := '0';
    --signal r_data_count : integer range 0 to OUTPUT_SIZE/8 := 0; -- Counter for received bytes

begin
    process(clk)
    begin
        if rising_edge(clk) then
            if i_DV = '1' then
                if r_status = '0' then
                    if r_input = r_condition then
                        r_status <= '1';
                    else
                        r_status <='0';                        
                    end if;
                end if;
            end if;
        end if;
    end process;
    o_status <= r_status;
    r_input <= i_input;
end behav;